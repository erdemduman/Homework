module xor_process(out, inA, inB);

input inA, inB;
output out;

xor two_inp_xor(out, inA, inB);

endmodule