module and_process(out, inA, inB);

input inA, inB;
output out;

and two_inp_and(out, inA, inB);

endmodule