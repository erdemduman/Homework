module or_process(out, inA, inB);

input inA, inB;
output out;

or two_inp_or(out, inA, inB);

endmodule